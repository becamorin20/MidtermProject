`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/13/2018 12:49:31 PM
// Design Name: 
// Module Name: CS151_controller
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module CS151_controller(
    input [31:0] inst,
    output [3:0] ALUopsel,
    output MUXsel1,
    output Regwrite
    );
endmodule
